module xm23_cpu (SW, HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, HEX6, HEX7, LEDG, LEDG7, LEDR, LEDR16_17, KEY, CLOCK_50, GPIO, KB_IN_GPIO, KB_OUT_GPIO, SCR_IN_GPIO, SCR_OUT_GPIO, test_gpio, test_gpio2);
	input [17:0] SW;
	input [3:0] KEY;
	input CLOCK_50;
	input GPIO;
	output wire [5:0] LEDG;
	output wire [15:0] LEDR;
	output reg [1:0] LEDR16_17;
	output reg LEDG7;
	output wire [6:0] HEX0;
	output wire [6:0] HEX1;
	output wire [6:0] HEX2;
	output wire [6:0] HEX3;
	output wire [6:0] HEX4;
	output wire [6:0] HEX5;
	output wire [6:0] HEX6;
	output wire [6:0] HEX7;

	input [8:0] KB_IN_GPIO;
	output wire KB_OUT_GPIO;
	output wire [8:0] SCR_OUT_GPIO;
	input SCR_IN_GPIO;
	output reg test_gpio;
	output reg test_gpio2;

	
	// Guide for memory initialization: https://projectf.io/posts/initialize-memory-in-verilog/
	// Example for how to initialize memory: https://stackoverflow.com/questions/70151532/read-from-file-to-memory-in-verilog

	reg [15:0] reg_file [0:16];			// Declare the register file
	reg [15:0] instr_reg, mar, mdr, psw_in;
	reg [15:0] data_bus, addr_bus;
	reg [2:0] ctrl_reg;
	reg execution_type = 1'b0;
	reg [15:0] bkpnt;
	reg [15:0] extension = 16'hffff;


	//devmem
	reg [7:0] dev_mem [0:15];

	// initial begin
	// 	dev_mem[0] = 8'b00010000;
	// 	dev_mem[1] = 8'b00000000;
	// 	dev_mem[2] = 8'b00010100;
	// 	dev_mem[3] = 8'b01101011;
	// 	dev_mem[4] = 8'b00000000;
	// 	dev_mem[5] = 8'b00000000;
	// end
	initial begin
		$readmemh("device_memory.txt", dev_mem, 0);
	end
	reg access_dev_mem;
	reg register_access_flag;
	reg word_rf_mdr;
	reg byte_rf_mdr;
	reg mar_not_used;
	wire [7:0] kb_data_output;
	parameter kb_csr = 0;
	parameter kb_data = 1;
	parameter scr_csr = 2;
	parameter scr_data = 3;
	parameter tmr_csr = 4;
	parameter tmr_data = 5;

	wire [7:0] arduino_data_i, arduino_data_o, csr_kb_o, csr_scr_o;
	wire [1:0] arduino_ctrl_i, arduino_ctrl_o;

	assign arduino_data_i = KB_IN_GPIO[7:0];
	assign arduino_data_o = SCR_OUT_GPIO[7:0];
	assign arduino_ctrl_o = {SCR_OUT_GPIO[8], KB_OUT_GPIO}; 
	assign arduino_ctrl_i = {KB_IN_GPIO[8], SCR_IN_GPIO};

	
	initial begin
		reg_file[0] = 16'd0;
		reg_file[1] = 16'd0;
		reg_file[2] = 16'd0;
		reg_file[3] = 16'd0;
		reg_file[4] = 16'd0;
		reg_file[5] = 16'd0;
		reg_file[6] = 16'h0800;
		reg_file[7] = 16'h1000;
		reg_file[8] = 16'd0;
		reg_file[9] = 16'd1;
		reg_file[10] = 16'd2;
		reg_file[11] = 16'd4;
		reg_file[12] = 16'd8;
		reg_file[13] = 16'd16;
		reg_file[14] = 16'd32;
		reg_file[15] = 16'hffff;
		reg_file[16] = 16'h0000;
		ctrl_reg = 3'b000;
		bkpnt = 16'h00f2;
		psw_in = 16'h60e0;
		mar = 16'h0000;
		mdr = 16'h0000;	
		
		register_access_flag = 1'b0;
	end
	
	wire Clock;
	wire [6:0] data_bus_ctrl, addr_bus_ctrl; 	// [1b for W/B, 3b for src, 3b for dst (Codes: 0=MDR/MAR, 1=Reg File, 2=IR, 3=ALU, 4=SXT_out, 5=BMB_out, 6=PSW)]
	wire s_bus_ctrl, sxt_bus_ctrl;							// 0 = use Reg File, 1 = use calculated offset
	wire [15:0] addr, breakpnt, PC;
	wire [4:0] dbus_rnum_dst, dbus_rnum_src, addr_rnum_src, alu_rnum_dst, alu_rnum_src, bm_rnum, sxt_rnum;
	wire [3:0] sxt_bit_num;
	wire [1:0] psw_bus_ctrl;
	wire [1:0] mem_mode;
	wire [15:0] mem_data, reg_data, psw_data;
	wire [15:0] mar_mem_bus, mdr_mem_bus;
	wire [15:0] sxt_in, sxt_out, alu_psw_out, psw_out;
	wire [15:0] bm_in, bm_out;
	wire [2:0] bm_op;
	wire [5:0] alu_op;
	wire [15:0] s_bus, d_bus, alu_out;
	wire [2:0] CR_bus;
	wire [3:0] cu_out1, cu_out2, cu_out3;
	wire id_E, ID_en;
	wire sxt_shift;
	
	wire [15:0] mem_ub_addr, mem_lb_addr;
	wire [7:0] mem_ub, mem_lb;
	
	wire [15:0] Instr;
	wire [6:0] OP;
	wire [12:0] OFF;
	wire [3:0] C;
	wire [2:0] T;
	wire [2:0] F;
	wire [2:0] PR;
	wire [3:0] SA;
	wire [4:0] PSWb;
	wire [2:0] DST;
	wire [2:0] SRCCON;
	wire WB;
	wire RC;
	wire [7:0] ImByte;
	wire PRPO;
	wire DEC;
	wire INC;
	wire ID_FLTo;
	wire [3:0] vect_num;
	wire [7:0] cex_state_out, cex_state_in;
	wire [1:0] PSW_ENT;
	wire pic_read, breakpnt_set;
	wire [7:0] pic_in;
	
	wire psw_update;
	wire [2:0] new_curr_pri;	// Priority of the new interrupt
	
	wire [3:0] nib4, nib5, nib6, nib7;
	
	assign pic_in = 8'b00000000;
	assign addr = SW[15:0];
	assign breakpnt = bkpnt[15:0];
	assign PC = reg_file[7][15:0];
	assign cex_state_in = mdr[7:0];
	
	assign mem_mode[1:0] = KEY[2:1];
	
	assign mem_data = mdr[15:0];
	assign psw_data = psw_out[15:0];
	assign reg_data = reg_file[addr[3:0]][15:0];
	
	//assign Clock = (execution_type == 1'b0) ? KEY[0] : CLOCK_50;
	assign Clock = GPIO;
	assign mar_mem_bus = mar[15:0];
	assign mem_ub_addr = (breakpnt_set == 1'b0) ? (mar[15:0] + 1) : (addr + 1);
	assign mem_lb_addr = (breakpnt_set == 1'b0) ? mar[15:0] : addr;
	
	assign new_curr_pri = reg_file[16][7:5];	// The new PSW is stored in the temp register (new pri accessed through this)
	
	assign d_bus = reg_file[alu_rnum_dst[4:0]][15:0];
	assign bm_in = reg_file[bm_rnum[3:0]][15:0];
	assign sxt_in = (sxt_bus_ctrl == 1'b0) ? reg_file[sxt_rnum[3:0]][15:0] : OFF[12:0];
	assign s_bus = (s_bus_ctrl == 1'b0) ? reg_file[alu_rnum_src[4:0]][15:0] : sxt_out[15:0];
	
	// Assign enable
	assign id_E = ID_en;
	
	assign nib4 = cu_out2[3:0];
	assign nib5 = cu_out3[3:0];
	assign nib6 = s_bus[3:0];
	assign nib7 = cu_out1;
	
	seven_seg_decoder decode5( .Reg1 (nib4), .HEX0 (HEX4), .Clock (Clock));
	seven_seg_decoder decode6( .Reg1 (nib5), .HEX0 (HEX5), .Clock (Clock));
	seven_seg_decoder decode7( .Reg1 (nib6), .HEX0 (HEX6), .Clock (Clock));
	seven_seg_decoder decode8( .Reg1 (nib7), .HEX0 (HEX7), .Clock (~Clock));
	
	
	memory ram(Clock, mdr[7:0], mdr[15:8], mem_lb_addr, mem_ub_addr, ctrl_reg[0], ctrl_reg[1], mem_lb, mem_ub);

	view_data data_viewer(mem_data, reg_data, psw_data, addr, KEY[3], mem_mode, HEX0, HEX1, HEX2, HEX3, LEDG, LEDR);
	
	sign_extender sxt_ext(sxt_in, sxt_out, sxt_bit_num, sxt_shift);
	
	byte_manip byte_manipulator(bm_op, bm_in, bm_out, ImByte);
	
	instruction_decoder ID(instr_reg, id_E, OP, OFF, C, T, F, PR, SA, PSWb, DST, SRCCON, WB, RC, ImByte, PRPO, DEC, INC, ID_FLTo, Clock);
	
	control_unit ctrl_unit(Clock, ID_FLTo, OP, OFF, C, T, F, PR, SA, PSWb, DST, SRCCON, WB, RC, PRPO, DEC, INC, psw_in, psw_out, 
							ID_en, CR_bus, data_bus_ctrl, addr_bus_ctrl, s_bus_ctrl, sxt_bit_num, sxt_rnum, sxt_shift, alu_op, 
							psw_update, dbus_rnum_dst, dbus_rnum_src, alu_rnum_dst, alu_rnum_src, sxt_bus_ctrl, bm_rnum, bm_op,
							breakpnt, PC, addr_rnum_src, psw_bus_ctrl, cu_out1, cu_out2, cu_out3, vect_num, PSW_ENT, cex_state_out,
							cex_state_in, new_curr_pri, pic_in, pic_read, breakpnt_set);
	
	alu arithmetic_logic_unit(d_bus, s_bus, alu_out, alu_op, psw_out, alu_psw_out, psw_update);

	kb_scr_drv kb_scr(	kb_data_output, dev_mem[scr_data][7:0], dev_mem[kb_csr][7:0], dev_mem[scr_csr][7:0], arduino_data_i, 
						arduino_data_o, arduino_ctrl_i, arduino_ctrl_o, csr_scr_o, csr_kb_o, Clock);

	// Indicator of whether CPU is currently executing instructions based on PSW SLP bit
	always @(psw_data[3]) begin
		if (psw_data[3] == 1'b1)
			LEDR16_17[0] = 1'b0;	// Not executing
		else
			LEDR16_17[0] = 1'b1;	// Executing
	end
	
	// Selection of execution modes. SW16 = 1 for continuous. SW16 = 0 for step.
	always @(SW[16]) begin
		if (SW[16] == 1'b1) begin
			LEDR16_17[1] = 1'b1;
			execution_type = 1'b1;
		end
		else begin
			LEDR16_17[1] = 1'b0;
			execution_type = 1'b0;
		end
	end
	
	// Breakpoint setting
	always @(SW[17]) begin
		if (SW[17] == 1'b1) begin
			LEDG7 = 1'b1;
			bkpnt <= addr[15:0];
		end
		else
			LEDG7 = 1'b0;
	end
	
	// Update registers
	always @(negedge Clock) begin
		ctrl_reg = CR_bus[2:0];
		if (psw_bus_ctrl == 2'b00)
			psw_in <= alu_psw_out[15:0];
		else if (psw_bus_ctrl == 2'b01)
			psw_in <= mdr[15:0];
		else if (psw_bus_ctrl == 2'b10)
			psw_in <= reg_file[dbus_rnum_src[4:0]][15:0];
		else if (psw_bus_ctrl == 2'b11)
			psw_in <= psw_data[15:0];
	end

	// Bus Assignment (MUX)
	always @(negedge Clock) begin
		access_dev_mem = 1'b0;
		register_access_flag = 1'b0;
		word_rf_mdr = 1'b0;
		byte_rf_mdr = 1'b0;
		mar_not_used = 1'b0;
		//clear flag
		
		//Address Bus Updating
		if (addr_bus_ctrl[2:0] == 3'b000) begin 			// MAR
			if (addr_bus_ctrl[5:3] == 3'b001)				// Read from Register File into MAR
				mar = reg_file[addr_rnum_src[4:0]][15:0];
			else if (addr_bus_ctrl[5:3] == 3'b011) 			// Read from ALU Output into MAR
				mar = alu_out[15:0];
			else if (addr_bus_ctrl[5:3] == 3'b100)			// Read from Interrupt Vector addresses
				mar = 16'hffc0 + (vect_num[3:0] << 2) + PSW_ENT[1:0];	// Determine address from vector number and option
		end	
		else if (addr_bus_ctrl[2:0] == 3'b111) begin
			mar_not_used = 1'b1;
		end

		if (mar <=16 && mar >=0) begin
			access_dev_mem = 1'b1;
		end

		
		mdr[7:0] = mem_lb[7:0];
		mdr[15:8] = mem_ub[7:0];
		
		// Data Bus Updating
		if (data_bus_ctrl[2:0] == 3'b000) begin 			// MDR
			if (data_bus_ctrl[5:3] == 3'b001) begin			// Read from Register File into MDR
				mdr = reg_file[dbus_rnum_src[4:0]][15:0]; 
				if(access_dev_mem) begin
					register_access_flag = 1'b1;
				end
			end
			else if (data_bus_ctrl[5:3] == 3'b011)			// Read from ALU Output into MDR
				mdr = alu_out[15:0];
			else if (data_bus_ctrl[5:3] == 3'b100)			// Read from PSW into MDR
				mdr = psw_data[15:0];
			else if (data_bus_ctrl[5:3] == 3'b101)			// Read from CEX into MDR
				mdr = 16'h0 + cex_state_out[7:0];
			// if (access_dev_mem) begin
				//dev_mem[mar[3:0]] = (!flag ? driver_output : mdr) ;
				//byte/word functionality
			// end
		end
		else if (data_bus_ctrl[2:0] == 3'b001) begin 		// Register File
			if (data_bus_ctrl[5:3] == 3'b000)				// Read from MDR into Register File
				if (data_bus_ctrl[6] == 1'b1)				// Byte
					reg_file[dbus_rnum_dst[4:0]][7:0] = mdr[7:0];
					if(access_dev_mem) begin
						byte_rf_mdr = 1'b1;
					end
				else										// Word
					reg_file[dbus_rnum_dst[4:0]] = mdr[15:0];
					if(access_dev_mem) begin
						word_rf_mdr = 1'b1;
					end
			else if (data_bus_ctrl[5:3] == 3'b011) begin	// Read from ALU Output into Register File
				if (data_bus_ctrl[6] == 1'b1)				// Byte
					reg_file[dbus_rnum_dst[4:0]][7:0] = alu_out[7:0];
				else										// Word
					reg_file[dbus_rnum_dst[4:0]] = alu_out[15:0];
			end
			else if (data_bus_ctrl[5:3] == 3'b001) begin 	// Read from Register File into Register File
				if (data_bus_ctrl[6] == 1'b1)				// Byte
					reg_file[dbus_rnum_dst[4:0]][7:0] = reg_file[dbus_rnum_src[4:0]][7:0];
				else										// Word
					reg_file[dbus_rnum_dst[4:0]] = reg_file[dbus_rnum_src[4:0]][15:0];
			end
			else if (data_bus_ctrl[5:3] == 3'b100) begin 	// Read from Sign Extender Output into Register File
				reg_file[dbus_rnum_dst[4:0]] = sxt_out[15:0];
			end
			else if (data_bus_ctrl[5:3] == 3'b101) begin 	// Read from Byte Manipulator Output into Register File
				reg_file[dbus_rnum_dst[4:0]] = bm_out[15:0];
			end
		end
		else if (data_bus_ctrl[2:0] == 3'b010) begin 		// Instruction Register
			if (data_bus_ctrl[5:3] == 3'b001)				// Read from Register File into Instruction Register
				instr_reg = reg_file[dbus_rnum_src[4:0]][15:0];
			else if (data_bus_ctrl[5:3] == 3'b000)			// Read from MDR into Instruction Register
				instr_reg = mdr[15:0];
		end
		
		dev_mem[kb_csr] = (!register_access_flag ? csr_kb_o : (mar[3:0] == kb_csr) ? mdr : dev_mem[kb_csr]);
		dev_mem[scr_csr] = (!register_access_flag ? csr_scr_o : (mar[3:0] == scr_csr) ? mdr : dev_mem[scr_csr]); //of/dba set here?
		if (register_access_flag && mar[3:0] == scr_data) begin
			dev_mem[scr_data] = mdr;
			if (~dev_mem[scr_csr][2]) begin //check dba
				dev_mem[scr_csr][3] = 1'b1;
			end
			dev_mem[scr_csr][2] = 1'b0;
		end
		dev_mem[kb_data][7:0] = kb_data_output;

		//read
		if(addr_bus_ctrl[2:0] != 3'b111) begin
			if (byte_rf_mdr) begin
				mdr = dev_mem[mar[3:0]][7:0];
			end
			else if (word_rf_mdr) begin
				mdr = dev_mem[mar[3:0]][7:0] << 8 | dev_mem[mar[3:0] + 1][7:0];
			end
		end
		if (byte_rf_mdr || word_rf_mdr) begin
				if(mar[3:0] == kb_csr) begin
					dev_mem[kb_csr][2] = 1'b0;//dev_mem[kb_csr] & ~(1'b1 << 2); //dba clear
					dev_mem[kb_csr][3] = 1'b0;//dev_mem[kb_csr] & ~(1'b1 << 3); //of clear
				end
			end
		//write
		//if register_access_flag
		// if(data_bus_ctrl == 7'b0001000) begin
		// 	if (mar == scr_data) begin
		// 	end

		// end

			// else if (mar[3:0] == scr_data) begin
			// 	dev_mem[scr_csr] = dev_mem[scr_csr] | 1'b1 << 2; //dba set
			// 	dev_mem[scr_csr] = dev_mem[scr_csr] & 1'b1 << 3; //of clear
			// end


			// dev_mem[tmr_csr] = (!register_access_flag ? driver_output_tmr : mdr);
			// dev_mem[tmr_data] = (!register_access_flag ? driver_output_tmr : mdr);

/*
			(!flag_2 ? drv_output : mdr) = devmem
			mdr = (!flag ? driver_output_kb : devmem[kb_csr]);
			mdr = (!flag ? driver_output_kb : devmem[kb_data]);
			mdr = (!flag ? driver_output_kb : devmem[scr_csr]);
			mdr = (!flag ? driver_output_kb : devmem[tmr_csr]);
		*/



	end
endmodule